module top(
    input sys_clk,
    input sys_rst_n
    );

    wire locked;
    wire reset = ~sys_rst_n || ~locked;
    
    // ===========================================================
    wire [31:0] PC, Instr, MemAddr, WriteData, ReadData;
    wire [3:0] MemWrite_EN;

    processor_core cpu (
        .clk (clk_core),
        .reset (reset),

        .PC (PC),
        .Instr (Instr),

        .MemWrite_EN (MemWrite_EN),
        .MemAddr (MemAddr),
        .WriteData (WriteData),
        .ReadData (ReadData)
    );

    clk_wiz_0 clk_wiz (
        .clk_in1 (sys_clk),
        .reset (~sys_rst_n),
        .locked (locked),
        .clk_out1 (clk_core)
    );

    INSTR_MEM imem (
        .clka (clk_core),
        .ena (1'b1),
        .wea (1'b0),    // instr read only
        .addra (PC[11:2]),
        .dina (32'b0),
        .douta (Instr)
    );

    // DMEM
    DATA_MEM dmem (
        .clka (clk_core),
        .ena (1'b1),
        .wea (MemWrite_EN),
        .addra (MemAddr[11:2]),
        .dina (WriteData),
        .douta (ReadData)
    );

endmodule
